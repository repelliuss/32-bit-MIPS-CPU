`define DELAY 20
module alu1_testbench();
   reg a, b, ci;
   reg [2:0] alu_code;
   reg exp_ri, exp_cip1;
   wire tresult;
   wire ri, cip1;

   alu1 al0(ri, cip1, a, b, ci, alu_code);

   wire t0, t1;
   xnor xn0(t0, ri, exp_ri);
   xnor xn1(t1, cip1, exp_cip1);
   and a0(tresult, t0, t1);

   initial begin
      a = 1'b1;
      b = 1'b0;
      ci= 1'b0;
      alu_code = 3'b000;
      exp_ri = 1'b0;
      exp_cip1 = 1'b0;
      #`DELAY;
      a = 1'b1;
      b = 1'b1;
      ci= 1'b0;
      alu_code = 3'b000;
      exp_ri = 1'b1;
      exp_cip1 = 1'b1;
      #`DELAY;
      a = 1'b1;
      b = 1'b0;
      ci= 1'b0;
      alu_code = 3'b001;
      exp_ri = 1'b1;
      exp_cip1 = 1'b0;
      #`DELAY;
      a = 1'b1;
      b = 1'b1;
      ci= 1'b0;
      alu_code = 3'b001;
      exp_ri = 1'b1;
      exp_cip1 = 1'b1;
      #`DELAY;
      a = 1'b0;
      b = 1'b0;
      ci= 1'b0;
      alu_code = 3'b001;
      exp_ri = 1'b0;
      exp_cip1 = 1'b0;
      #`DELAY;
      a = 1'b0;
      b = 1'b0;
      ci= 1'b0;
      alu_code = 3'b010;
      exp_ri = 1'b0;
      exp_cip1 = 1'b0;
      #`DELAY;
      a = 1'b0;
      b = 1'b1;
      ci= 1'b0;
      alu_code = 3'b010;
      exp_ri = 1'b1;
      exp_cip1 = 1'b0;
      #`DELAY;
      a = 1'b1;
      b = 1'b1;
      ci= 1'b0;
      alu_code = 3'b010;
      exp_ri = 1'b0;
      exp_cip1 = 1'b1;
      #`DELAY;
      a = 1'b1;
      b = 1'b1;
      ci= 1'b1;
      alu_code = 3'b010;
      exp_ri = 1'b1;
      exp_cip1 = 1'b1;
      #`DELAY;
      a = 1'b1;
      b = 1'b1;
      ci= 1'b1;
      alu_code = 3'b110;
      exp_ri = 1'b0;
      exp_cip1 = 1'b1;
      #`DELAY;
      a = 1'b1;
      b = 1'b0;
      ci= 1'b1;
      alu_code = 3'b110;
      exp_ri = 1'b1;
      exp_cip1 = 1'b1;
      #`DELAY;
      a = 1'b0;
      b = 1'b0;
      ci= 1'b1;
      alu_code = 3'b110;
      exp_ri = 1'b0;
      exp_cip1 = 1'b1;
      #`DELAY;
      a = 1'b1;
      b = 1'b1;
      ci= 1'b0;
      alu_code = 3'b011;
      exp_ri = 1'b0;
      exp_cip1 = 1'b1;
      #`DELAY;
      a = 1'b1;
      b = 1'b0;
      ci= 1'b0;
      alu_code = 3'b011;
      exp_ri = 1'b1;
      exp_cip1 = 1'b0;
      #`DELAY;
      a = 1'b0;
      b = 1'b1;
      ci= 1'b0;
      alu_code = 3'b011;
      exp_ri = 1'b1;
      exp_cip1 = 1'b0;
      #`DELAY;
      a = 1'b0;
      b = 1'b0;
      ci= 1'b0;
      alu_code = 3'b011;
      exp_ri = 1'b0;
      exp_cip1 = 1'b0;
   end

   initial begin
      $monitor("time = %2d, a =%1b, b=%1b, ci=%1b,  alu_code=%3b, ri=%1b, exp_ri=%1b, cip1=%1b, exp_cip1=%1b, tresult=%1b", $time, a, b, ci,alu_code, ri, exp_ri, cip1, exp_cip1, tresult);
   end

endmodule //alu1_testbench
